library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use work.types.all;

---------------------------------------------- ***** Description ***** ----------------------------------------------
-- Returns the absolute positions of each piece of the requested tile
-- This module is used to:
--	- * Write movements *
-- - * Check overlapping *
---------------------------------------------------------------------------------------------------------------------

entity tiles_memory is
	port (----------------
			---- INPUTS ----
			----------------
			tile		: in STD_LOGIC_VECTOR(5-1 downto 0);
			rotation : in STD_LOGIC_VECTOR(3-1 downto 0);			
			-----------------
			---- OUTPUTS ----
			-----------------
			tile_definition: out STD_LOGIC_VECTOR(102-1 downto 0)
	);
end tiles_memory;

architecture tiles_memoryArch of tiles_memory is
	-- Tiles memory
	-- ROM
	type ROM_type is array(0 to 168-1) of STD_LOGIC_VECTOR(102-1 downto 0);
	signal ROM: ROM_type :=(-- U
									"000101000001101000001000000000111111111111111111111111101101110000101001000110001101000010001001010000",
									"000101000001101000001000000000111111111111111111111111101101110000101001000110001101000010001001010000",
									"000101000001101000001000000000111111111111111111111111101101110000101001000110001101000010001001010000",
									"000101000001101000001000000000111111111111111111111111101101110000101001000110001101000010001001010000",
									"000101000001101000001000000000111111111111111111111111101101110000101001000110001101000010001001010000",
									"000101000001101000001000000000111111111111111111111111101101110000101001000110001101000010001001010000",
									"000101000001101000001000000000111111111111111111111111101101110000101001000110001101000010001001010000",
									"000101000001101000001000000000111111111111111111111111101101110000101001000110001101000010001001010000",
									-- T
									"000001001000101000101101000000111111111111111111101110110101000101110000101001000010001001001101010000",
									"000001001000101000001101000000111111111111111111101101110000101001000101000010001001001110010101010000",
									"000001101000001101000101000000111111111111111111101101110000101001000110001000000010001001001110010101",
									"000001001000000101101101000000111111111111111111101110110101101000000110001101101001000010001001010000",
									"001001001000101000000101000000111111111111111111101101110000101001000110001101000001010000001010010001",
									"101001001000101000000101000000111111111111111111101101110000110001101010000001000110001101001001010000",
									"000001101001001000000101000000111111111111111111101000110001101010000110101101001101000010001001010000",
									"001001000001101000000101000000111111111111111111101101110000101001000110001101001000000010001010010001",
									-- S
									"001001001000101000101101000000111111111111101110110101000101110000101001000001001101010000001010010001",
									"101001001000101000001101000000111111111111101101110000110001101010000001000101001110010101001001010000",
									"000001101001001101000101000000111111111111101000110001101010000110101101001000000010001001001110010101",
									"001001000001000101101101000000111111111111101110110101101000000110001101001000101001000010001010010001",
									"001001001000101000101101000000111111111111101110110101000101110000101001000001001101010000001010010001",
									"101001001000101000001101000000111111111111101101110000110001101010000001000101001110010101001001010000",
									"000001101001001101000101000000111111111111101000110001101010000110101101001000000010001001001110010101",
									"001001000001000101101101000000111111111111101110110101101000000110001101001000101001000010001010010001",
									-- R
									"001001001000000101101101000000111111111111111111101110110101101000000110001101000001010000001010010001",
									"101001101000001101000101000000111111111111111111101101110000110001101010000001000110001000001110010101",
									"000001101001001000001101000000111111111111111111101000110001101010000101000010001001001110010101010000",
									"001001000001101000101101000000111111111111111111101110110101000101110000101001001000000010001010010001",
									"001001000001101000101101000000111111111111111111101110110101000101110000101001001000000010001010010001",
									"000001101001001000001101000000111111111111111111101000110001101010000101000010001001001110010101010000",
									"101001101000001101000101000000111111111111111111101101110000110001101010000001000110001000001110010101",
									"001001001000000101101101000000111111111111111111101110110101101000000110001101000001010000001010010001",									
									-- Q
									"010000001000000101000110000000111111000111101110001110101101001101101000000001001001010101010001011000",
									"110000101000000101000110000000111111110101111000110001101101101001000111101110001110001101000001001000",
									"010000001000000001000010000000111111000101101000101001001001101010000011001010001101010101010001011000",
									"110000101000000001000010000000111111110101111000110001101101101001000101001000001001101010000011001010",
									"110000101000000001000010000000111111110101111000110001101101101001000101001000001001101010000011001010",
									"010000001000000001000010000000111111000101101000101001001001101010000011001010001101010101010001011000",
									"110000101000000101000110000000111111110101111000110001101101101001000111101110001110001101000001001000",
									"010000001000000101000110000000111111000111101110001110101101001101101000000001001001010101010001011000",
									-- P
									"000101001001000001101001000000111111111111101000110001101010000110101101001101001000000010001010010001",
									"000101001001000001101001000000111111111111101000110001101010000110101101001101001000000010001010010001",
									"001000101001101000101101000000111111111111101110110101000101110000110001101010000001001101001001010000",
									"101000001001001000001101000000111111111111101101110000101001000101000001001110010101010000001010010001",
									"000001001101000101101101000000111111111111101110110101101000000110001000101001000010001001001110010101",
									"000001001101000101101101000000111111111111101110110101101000000110001000101001000010001001001110010101",
									"101000001001001000001101000000111111111111101101110000101001000101000001001110010101010000001010010001",
									"001000101001101000101101000000111111111111101110110101000101110000110001101010000001001101001001010000",
									-- O
									"001000000010000001000101000000111111111111000110101101001101101000101001001001101010000011001010010000",
									"101000000010000001000101000000111111111111101101110000101001000110001101001000001001101010000011001010",
									"000001110000101000001000000000111111111111110101111000110001101101101001000101000010001001001101010000",
									"000001010000001000101000000000111111111111101101110000101001000101000010001001001101010101010001011000",
									"101000000110000101000001000000111111111111101101110000101001000111101110001110001101001000000010001001",
									"001000000110000101000001000000111111111111000111101110001110101101001101101000101001000010001001010000",
									"000101010000001000101000000000111111111111101101110000101001000110001101000001001001010101010001011000",
									"000101110000101000001000000000111111111111110101111000110001101101101001000110001101000001001001010000",
									-- N
									"101001101101000001000101000000111111111111101110110101101000110001101010000110001101001000000010001001",
									"001101001001000001000101000000111111111111000110101101101000001000101001000010001110010101001010010001",
									"101101001101001000101000000000111111111111101110110101000101110000101001000001001110010101001001010000",
									"101101001101001000101000000000111111111111101110110101000101110000101001000001001110010101001001010000",
									"001101001001000001000101000000111111111111000110101101101000001000101001000010001110010101001010010001",
									"101001101101000001000101000000111111111111101110110101101000110001101010000110001101001000000010001001",
									"001001101001001000101000000000111111111111101101110000110001101010000001000101001101010000001010010001",
									"001001101001001000101000000000111111111111101101110000110001101010000001000101001101010000001010010001",
									-- M
									"101001101000000001000101000000111111111111111111101101110000110001101010000110001101001000000010001001",
									"001001001000000001000101000000111111111111111111000110101101001101101000101001000010010000001010010001",
									"101101000101001000101000000000111111111111111111101110110101110000101001000110001101000001001001010000",
									"001101000101001000101000000000111111111111111111101101110000101001000110000001001110010101001001010000",
									"001101001000000001000101000000111111111111111111000110101101101000101001000010001001001110010101010000",
									"101101101000000001000101000000111111111111111111101110110101110000101001000110001101001000000010001001",
									"001001000001001000101000000000111111111111111111101101110000101001000101000010001101010000001010010001",
									"101001000001001000101000000000111111111111111111101101110000110001101010000101000010001001001101010000",
									-- L
									"101001101000000110000101000000111111111111101101110000110001101010000001000111101110001110001101001000",
									"001001001000000110000101000000111111111111000111101110001110101101001101101000000001010000001010010001",
									"101101000101010000001000000000111111111111101110110101101000000110001101000001001001010101010001011000",
									"001101000101110000101000000000111111111111110101111000110001101101101001000110000001001000001110010101",
									"001101001000000010000001000000111111111111000101101000101001001001101010000011001010001110010101010000",
									"101101101000000010000001000000111111111111101110110101000101110000101001001000001001101010000011001010",
									"001001000001110000101000000000111111111111110101111000110001101101101001000101001000000010001010010001",
									"101001000001010000001000000000111111111111101000110001101010000101000010001001001101010101010001011000",
									-- K
									"101001000001000101000110000000111111101000110001101010000111101110001110101101001101001000000010001001",
									"001001000001000101000110000000111111000111101110001110101101001101101000001000101001000010001010010001",
									"101101010000001000101000000000111111101110110101000101110000101001000001001101001001010101010001011000",
									"001101001000101000110000000000111111110101111000110001101101101001000101000001001110010101001001010000",
									"001101000010000001000101000000111111000110101101101000001000101001001001101010000011001010001110010101",
									"101101000010000001000101000000111111101110110101101000000110001101001000101001001001101010000011001010",
									"001001001000101000110000000000111111110101111000110001101101101001000101000001001101010000001010010001",
									"101001010000001000101000000000111111101101110000110001101010000001000101001101001001010101010001011000",
									-- J
									"000110000101000010000001000000000111101110001110101101001101101000001000101001001001101010000011001010",
									"000110000101000010000001000000000111101110001110101101001101101000001000101001001001101010000011001010",
									"110000101000010000001000000000110101111000110001101101101001000101000001001101001001010101010001011000",
									"110000101000010000001000000000110101111000110001101101101001000101000001001101001001010101010001011000",
									"000110000101000010000001000000000111101110001110101101001101101000001000101001001001101010000011001010",
									"000110000101000010000001000000000111101110001110101101001101101000001000101001001001101010000011001010",
									"110000101000010000001000000000110101111000110001101101101001000101000001001101001001010101010001011000",
									"110000101000010000001000000000110101111000110001101101101001000101000001001101001001010101010001011000",									
									-- I
									"111111001001000001101000000000111111111111111111111111101101110000101001000101001000000010001010010001",
									"111111101001000001001000000000111111111111111111111111101000110001101010000101000010001001001101010000",
									"111111000101101001101000000000111111111111111111111111101101110000110001101010000001000110001101001000",
									"111111000101001001001000000000111111111111111111111111000110101101001101101000000001010000001010010001",
									"111111101101000101001000000000111111111111111111111111101110110101101000000110001101000001001001010000",
									"111111001101000101101000000000111111111111111111111111101101110000101001000110000001001000001110010101",
									"111111001101000001001000000000111111111111111111111111000101101000101001000010001001001110010101010000",
									"111111101101000001101000000000111111111111111111111111101110110101000101110000101001001000000010001001",
									-- H
									"111111001001000001001000000000111111111111111111111111000101101000101001000010001101010000001010010001",
									"111111101001000001101000000000111111111111111111111111101101110000110001101010000101001000000010001001",
									"111111101001000001101000000000111111111111111111111111101101110000110001101010000101001000000010001001",
									"111111001001000001001000000000111111111111111111111111000101101000101001000010001101010000001010010001",
									"111111101101000101101000000000111111111111111111111111101110110101110000101001000110001101000001001000",
									"111111001101000101001000000000111111111111111111111111000110101101101000000001001110010101001001010000",
									"111111001101000101001000000000111111111111111111111111000110101101101000000001001110010101001001010000",
									"111111101101000101101000000000111111111111111111111111101110110101110000101001000110001101000001001000",
									-- G
									"111111001000000101000001000000111111111111111111111111000110101101001101101000101001000010001001010000",
									"111111101000000101000001000000111111111111111111111111101101110000101001000110001101001000000010001001",
									"111111000001101000001000000000111111111111111111111111101101110000101001000101000010001001001101010000",
									"111111000001101000001000000000111111111111111111111111101101110000101001000101000010001001001101010000",
									"111111101000000101000001000000111111111111111111111111101101110000101001000110001101001000000010001001",
									"111111001000000101000001000000111111111111111111111111000110101101001101101000101001000010001001010000",
									"111111000101101000001000000000111111111111111111111111101101110000101001000110001101000001001001010000",
									"111111000101101000001000000000111111111111111111111111101101110000101001000110001101000001001001010000",
									-- F
									"111111101001000001000101000000111111111111111111101000110001101010000110101101001101001000000010001001",
									"111111001001000001000101000000111111111111111111000110101101001101101000001000101001000010001010010001",
									"111111101101101000001000000000111111111111111111101110110101000101110000101001000001001101001001010000",
									"111111001101101000001000000000111111111111111111101101110000101001000101000001001110010101001001010000",
									"111111001101000101000001000000111111111111111111000110101101101000001000101001000010001001001110010101",
									"111111101101000101000001000000111111111111111111101110110101101000000110001101001000101001000010001001",
									"111111001001101000001000000000111111111111111111101101110000101001000101000001001101010000001010010001",
									"111111101001101000001000000000111111111111111111101101110000110001101010000001000101001101001001010000",
									-- E
									"111111000010000001000101000000111111111111000110101101001101101000001000101001001001101010000011001010",
									"111111000010000001000101000000111111111111000110101101001101101000001000101001001001101010000011001010",
									"111111001000110000101000000000111111111111110101111000110001101101101001000101000001001101001001010000",
									"111111010000001000101000000000111111111111101101110000101001000101000001001101001001010101010001011000",
									"111111000110000101000001000000111111111111000111101110001110101101001101101000001000101001000010001001",
									"111111000110000101000001000000111111111111000111101110001110101101001101101000001000101001000010001001",
									"111111010000001000101000000000111111111111101101110000101001000101000001001101001001010101010001011000",
									"111111001000110000101000000000111111111111110101111000110001101101101001000101000001001101001001010000",
									-- D
									"111111111111000101001000000000111111111111111111111111111111000110101101001101101000000001001001010000",
									"111111111111000101101000000000111111111111111111111111111111101101110000101001000110001101000001001000",
									"111111111111000001001000000000111111111111111111111111111111000101101000101001000010001001001101010000",
									"111111111111101000000001000000111111111111111111111111111111101101110000101001000101001000000010001001",
									"111111111111101000000001000000111111111111111111111111111111101101110000101001000101001000000010001001",
									"111111111111000001001000000000111111111111111111111111111111000101101000101001000010001001001101010000",
									"111111111111000101101000000000111111111111111111111111111111101101110000101001000110001101000001001000",
									"111111111111000101001000000000111111111111111111111111111111000110101101001101101000000001001001010000",
									-- C
									"111111111111000101000001000000111111111111111111111111000110101101001101101000001000101001000010001001",
									"111111111111000101000001000000111111111111111111111111000110101101001101101000001000101001000010001001",
									"111111111111101000001000000000111111111111111111111111101101110000101001000101000001001101001001010000",
									"111111111111101000001000000000111111111111111111111111101101110000101001000101000001001101001001010000",
									"111111111111000101000001000000111111111111111111111111000110101101001101101000001000101001000010001001",
									"111111111111000101000001000000111111111111111111111111000110101101001101101000001000101001000010001001",
									"111111111111101000001000000000111111111111111111111111101101110000101001000101000001001101001001010000",
									"111111111111101000001000000000111111111111111111111111101101110000101001000101000001001101001001010000",
									-- B
									"111111111111111111000001000000111111111111111111111111111111111111000101101000001000101001000010001001",
									"111111111111111111000001000000111111111111111111111111111111111111000101101000001000101001000010001001",
									"111111111111111111101000000000111111111111111111111111111111111111101101110000101001000101000001001000",
									"111111111111111111001000000000111111111111111111111111111111111111000101101000000001001101001001010000",
									"111111111111111111000101000000111111111111111111111111111111111111000110101101001101101000000001001000",
									"111111111111111111000101000000111111111111111111111111111111111111000110101101001101101000000001001000",
									"111111111111111111001000000000111111111111111111111111111111111111000101101000000001001101001001010000",
									"111111111111111111101000000000111111111111111111111111111111111111101101110000101001000101000001001000",
									-- A
									"111111111111111111111111000000111111111111111111111111111111111111111111111111000101101000000001001000",
									"111111111111111111111111000000111111111111111111111111111111111111111111111111000101101000000001001000",
									"111111111111111111111111000000111111111111111111111111111111111111111111111111000101101000000001001000",
									"111111111111111111111111000000111111111111111111111111111111111111111111111111000101101000000001001000",
									"111111111111111111111111000000111111111111111111111111111111111111111111111111000101101000000001001000",
									"111111111111111111111111000000111111111111111111111111111111111111111111111111000101101000000001001000",
									"111111111111111111111111000000111111111111111111111111111111111111111111111111000101101000000001001000",
									"111111111111111111111111000000111111111111111111111111111111111111111111111111000101101000000001001000");

	signal tiles_mem_addr: STD_LOGIC_VECTOR(8-1 downto 0);
begin
	-- Address
	tiles_mem_addr <= tile & rotation;
	
	-- Output
	tile_definition <= ROM(conv_integer(tiles_mem_addr));
end tiles_memoryArch;